localparam ALU8_ADD = 3'b000;
localparam ALU8_ADC = 3'b001;
localparam ALU8_SUB = 3'b010;
localparam ALU8_SBC = 3'b011;
localparam ALU8_OR  = 3'b100;
localparam ALU8_AND = 3'b101;
localparam ALU8_XOR = 3'b110;
localparam ALU8_LD  = 3'b111;