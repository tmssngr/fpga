localparam STATES_MAX_BIT = 4;
localparam STATE_FETCH_INSTR  = 0;
localparam STATE_READ_INSTR   = 1;
localparam STATE_WAIT_2       = 2;
localparam STATE_READ_2       = 3;
localparam STATE_WAIT_3       = 4;
localparam STATE_READ_3       = 5;
localparam STATE_DECODE       = 6;
localparam STATE_ALU1_WORD    = 7;
localparam STATE_ALU1_OP      = 8;
localparam STATE_ALU1_DA      = 9;
localparam STATE_ALU2_IR      = 10;
localparam STATE_ALU2_OP      = 11;
localparam STATE_PUSH         = 12;
localparam STATE_POP          = 13;
localparam STATE_DJNZ1        = 14;
localparam STATE_DJNZ2        = 15;
localparam STATE_LDC_READ     = 16;
localparam STATE_LDC_WRITE1   = 17;
localparam STATE_LDC_WRITE2   = 18;
localparam STATE_READ_MEM1    = 19;
localparam STATE_READ_MEM2    = 20;
localparam STATE_WRITE_MEM    = 21;
