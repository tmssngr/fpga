// similar to the upper nibble of the commands
localparam ALU8_ADD = 4'b0000;
localparam ALU8_ADC = 4'b0001;
localparam ALU8_SUB = 4'b0010;
localparam ALU8_SBC = 4'b0011;
localparam ALU8_OR  = 4'b0100;
localparam ALU8_AND = 4'b0101;
localparam ALU8_TCM = 4'b0110;
localparam ALU8_TM  = 4'b0111;
// 8
// 9
localparam ALU8_CP  = 4'b1010;
localparam ALU8_XOR = 4'b1011;
// c
// d
// e
localparam ALU8_LD  = 4'b1111;