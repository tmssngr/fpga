localparam ALU8_ADD = 2'b00;
localparam ALU8_LD = 2'b10;